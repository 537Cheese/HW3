module DECODER3 (Din, en, Dout);
parameter N = 32;
input [4:0] Din;
input en;
output [N-1 : 0] Dout;

assign {Dout} = 
( {en,Din} == 6'b100000) ? 32'b00000000000000000000000000000001 : 

( {en,Din} == 6'b100001) ? 32'b00000000000000000000000000000010 : 

( {en,Din} == 6'b100010) ? 32'b00000000000000000000000000000100 : 

( {en,Din} == 6'b100011) ? 32'b00000000000000000000000000001000 : 

( {en,Din} == 6'b100100) ? 32'b00000000000000000000000000010000 : 

( {en,Din} == 6'b100101) ? 32'b00000000000000000000000000100000 : 

( {en,Din} == 6'b100110) ? 32'b00000000000000000000000001000000 : 

( {en,Din} == 6'b100111) ? 32'b00000000000000000000000010000000 :
 
( {en,Din} == 6'b101000) ? 32'b00000000000000000000000100000000 : 

( {en,Din} == 6'b101001) ? 32'b00000000000000000000001000000000 :

( {en,Din} == 6'b101010) ? 32'b00000000000000000000010000000000 :

( {en,Din} == 6'b101011) ? 32'b00000000000000000000100000000000 :   

( {en,Din} == 6'b101100) ? 32'b00000000000000000001000000000000 : 

( {en,Din} == 6'b101101) ? 32'b00000000000000000010000000000000 : 

( {en,Din} == 6'b101110) ? 32'b00000000000000000100000000000000 : 

( {en,Din} == 6'b101111) ? 32'b00000000000000001000000000000000 : 

( {en,Din} == 6'b110000) ? 32'b00000000000000010000000000000000 : 

( {en,Din} == 6'b110001) ? 32'b00000000000000100000000000000000 : 

( {en,Din} == 6'b110010) ? 32'b00000000000001000000000000000000 : 

( {en,Din} == 6'b110011) ? 32'b00000000000010000000000000000000 : 

( {en,Din} == 6'b110100) ? 32'b00000000000100000000000000000000 : 

( {en,Din} == 6'b110101) ? 32'b00000000001000000000000000000000 : 

( {en,Din} == 6'b110110) ? 32'b00000000010000000000000000000000 : 

( {en,Din} == 6'b110111) ? 32'b00000000100000000000000000000000 : 

( {en,Din} == 6'b111000) ? 32'b00000001000000000000000000000000 : 

( {en,Din} == 6'b111001) ? 32'b00000010000000000000000000000000 : 

( {en,Din} == 6'b111010) ? 32'b00000100000000000000000000000000 : 

( {en,Din} == 6'b111011) ? 32'b00001000000000000000000000000000 : 

( {en,Din} == 6'b111100) ? 32'b00010000000000000000000000000000 : 

( {en,Din} == 6'b111101) ? 32'b00100000000000000000000000000000 : 

( {en,Din} == 6'b111110) ? 32'b01000000000000000000000000000000 : 

( {en,Din} == 6'b111111) ? 32'b10000000000000000000000000000000 : 32'b11111111111111111111111111111111;

endmodule
