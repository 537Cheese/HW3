`timescale 1ns/1ps
module MUX_TESTBENCH;

	reg[7:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31;

	
	reg[4:0] s;
	wire [7:0] o;

	MUX3 dut (o, i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,i31, s);
	
	initial 
	s = 5'b00000;
	always begin
	# 10 s = s + 1'b1;
	end
	
	initial begin
		i0<=8'b00000001;
		i1<=8'b00000010;
		i2<=8'b00000100;
		i3<=8'b00001000;
		i4<=8'b00010000;
		i5<=8'b00100000;
		i6<=8'b01000000;
		i7<=8'b10000000;
		i8<=8'b00000001;
		i9<=8'b00000010;
		i10<=8'b00000100;
		i11<=8'b00001000;
		i12<=8'b00010000;
		i13<=8'b00100000;
		i14<=8'b01000000;
		i15<=8'b10000000;
		i16<=8'b00000001;
		i17<=8'b00000010;
		i18<=8'b00000100;
		i19<=8'b00001000;
		i20<=8'b00010000;
		i21<=8'b00100000;
		i22<=8'b01000000;
		i23<=8'b10000000;
		i24<=8'b00000001;
		i25<=8'b00000010;
		i26<=8'b00000100;
		i27<=8'b00001000;
		i28<=8'b00010000;
		i29<=8'b00100000;
		i30<=8'b01000000;
		i31<=8'b10000000;
	end

	initial begin 
	#500 $stop;
	end
endmodule
